// ******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.1 D filp-flop        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
//
module top_module (
    input clk,    // Clocks are used in sequential circuits
    input d,
    output reg q );//

    always @(posedge clk ) begin
    	q <= d;
    end

endmodule


// ******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.2 D filp-flops       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input [7:0] d,
    output [7:0] q
);
    always @(posedge clk ) begin
    	q <= d;
    end

endmodule

// ******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.3 DFF with reset     /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input reset,            // Synchronous reset
    input [7:0] d,
    output [7:0] q
);
  always @(posedge clk ) begin
      if (reset) begin
  		q <= 7'b0;
  	end else begin
  		q <= d;
  	
  	end
  end
endmodule


// **************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.4 DFF with reset value       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input reset,
    input [7:0] d,
    output [7:0] q
);
  always @(negedge clk ) begin
      if (reset) begin
  		q <= 7'h34;
  	end else begin
  		q <= d;

  	end
  end
endmodule


// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.5 DFF with asynchronous reset   /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
  input clk,
  input areset,   // active high asynchronous reset
  input [7:0] d,
  output [7:0] q
);
always @(posedge clk or posedge areset) begin
	if ( areset ) begin
		 q <= 7'b00;
	end else begin
		 q <= d;
	end
end

endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.6 DFF with byte enable          /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input resetn,
    input [1:0] byteena,
    input [15:0] d,
    output [15:0] q
);
  always @ (posedge clk) begin
  	if (!resetn) begin
  		q <= 15'b0;
  	end else begin
  		q[7: 0] <= (byteena[0]) ? d[7: 0] : q[7: 0];
  		q[15: 8] <= (byteena[1]) ? d[15: 8] : q[15: 8];
  	end
  end

endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.7 D Latch                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input d,
    input ena,
    output q);
  assign q = (ena) ? d : q;

endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.8 DFF                           /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input d,
    input ar,   // asynchronous reset
    output q
);
  always @(posedge clk or posedge ar) begin
  	if ( ar ) begin
  		 q <= 1'b0;
  	end else begin
  		 q <= d;

  	end
  end
endmodule


// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.9 DFF                           /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input d,
    input r,   // synchronous reset
    output q
  );
	always @ (posedge clk) begin
		if (r) begin
			q <= 1'b0;
		end else begin
			q <= d;

		end
	end
endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.10 DFF+gate                     /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input in,
    output out
  );
	always_ff @(posedge clk) begin
		out <= out ^ in;
	end

endmodule


// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.11 Mux and DFF                  /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
//Mt2015 muxdff
module top_module (
	input clk,
	input L,
	input r_in,
	input q_in,
	output reg Q
);
  always @ (posedge clk) begin
  	if (L) begin
  		Q <= r_in;
  	end else begin
  		Q <= q_in;


  	end
  end
endmodule


// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.12 Mux and DFF                  /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
// 寫法1
module top_module (
    input clk,
    input w, R, E, L,
    output Q
);
	always @ (posedge clk) begin
  	if (E) begin
  		Q <= (L) ? R : w ;
  	end else begin
  		Q <= (L) ? R : Q ;
  	end
  end

endmodule

// 寫法2
module top_module (
    input clk,
    input w, R, E, L,
    output Q
);
    always@(posedge clk)begin
        Q <= L ? R : (E ? w : Q);
    end

endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.13 DFFs and gates               /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input x,
    output z
);
  reg [2:0] q;
	always @ (posedge clk) begin
		q[0] <= x ^  q[0];
		q[1] <= x & !q[1];
		q[2] <= x | !q[2];
	end

	assign z = !(|q);

endmodule

// *********************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/*
// S03-2-1.14 Create circuit from truth table  /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**
// *******************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/
// JK FF
module top_module (
    input clk,
    input j,
    input k,
    output Q
);
	always @ (posedge clk) begin
		case({j,k})
			2'b00: Q <= Q;
			2'b01: Q <= 1'b0;
			2'b10: Q <= 1'b1;
			2'b11: Q <= ~Q;
		endcase
	end

endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.15 Detect an edge               /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input [7:0] in,
    output [7:0] pedge
);
	reg [7: 0]  in_d1;

	always @(posedge clk) begin
		in_d1 <= in;
		pedge <= ~in_d1 & in;
	end
endmodule

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.16 Detect both edges            /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
module top_module (
    input clk,
    input [7:0] in,
    output [7:0] anyedge
);
	reg [7: 0]  in_d1;

	always @(posedge clk) begin
		in_d1 <= in;
		anyedge <= (~in_d1 & in) | (in_d1 & ~in);
	end
endmodule


// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.17 Edge capture register        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ******************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
// S03-2-1.18 Dual-edge triggered flip-flop /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****



