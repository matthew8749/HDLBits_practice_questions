// *****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.1 Simple FSM 1 (asynchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_1.Simple_FSM_1_(asynchronous reset)   // 無意義，快速找題目用
module top_module(
    input clk,
    input areset,    // Asynchronous reset to state B
    input in,
    output out
);//
    parameter A=0;
    parameter B=1;
    reg state;
    reg next_state;
    reg st_out;

    always @(*) begin    // This is a combinational always block
        if (areset) begin
        	next_state = B;
        end else begin
        	case (state)
        	B:  next_state = (in) ? B : A;
        	A:  next_state = (in) ? A : B;
        	default : next_state = B;
          endcase

        end
    end


		always @(posedge clk or posedge areset) begin    // This is a sequential always block
        // State flip-flops with asynchronous reset
        if ( areset ) begin
        	state <= B;
        end else begin
        	state <= next_state;

        end
    end

    always @(posedge clk or posedge areset) begin    // This is a sequential always block
        // State flip-flops with asynchronous reset
        if ( areset ) begin
        	st_out <= 1;
        end else begin
        	case (next_state)
        	  A: st_out <= 1'b0;
        	  B: st_out <= 1'b1;
        		default : st_out <= 1'b1;
        	endcase

        end
    end

    // Output logic
    assign out = st_out;

endmodule

// ****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.2 Simple FSM 1 (synchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_2.Simple_FSM_1_(synchronous reset)   // 無意義，快速找題目用
module top_module(
    input clk,
    input reset,    // Asynchronous reset to state B
    input in,
    output out
);//
    parameter A=0;
    parameter B=1;
    reg state;
    reg next_state;
    reg st_out;

    always @(*) begin    // This is a combinational always block
        if (reset) begin
        	next_state = B;
        end else begin
        	case (state)
        	B:  next_state = (in) ? B : A;
        	A:  next_state = (in) ? A : B;
        	default : next_state = B;
          endcase

        end
    end


		always @(posedge clk) begin    // This is a sequential always block
        // State flip-flops with asynchronous reset
        if ( reset ) begin
        	state <= B;
        end else begin
        	state <= next_state;

        end
    end

    always @(posedge clk) begin    // This is a sequential always block
        // State flip-flops with asynchronous reset
        if ( reset ) begin
        	st_out <= 1;
        end else begin
        	case (next_state)
        	  A: st_out <= 1'b0;
        	  B: st_out <= 1'b1;
        		default : st_out <= 1'b1;
        	endcase

        end
    end

    // Output logic
    assign out = st_out;

endmodule
// *****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.3 Simple FSM 2 (asynchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_3.Simple_FSM_2_(asynchronous reset)   // 無意義，快速找題目用
module top_module(
  input clk,
  input areset,    // Asynchronous reset to OFF
  input j,
  input k,
  output out
);

	parameter st_OFF=0;
  parameter st_ON=1;
  reg state;
  reg next_state;

  always @ (*) begin
  	if ( areset ) begin
  		 next_state = 0;
  	end else begin
  		case (state)
      st_OFF : next_state = (j) ? st_ON : st_OFF;
      st_ON  : next_state = (k) ? st_OFF: st_ON;
      default: next_state = (j) ? st_ON : st_OFF;
  		endcase

  	end
  end

  always @(posedge clk or posedge areset) begin
  	if ( areset ) begin
  		state <= st_OFF;
  	end else begin
  		state <= next_state;
  	end
  end

  assign out = (state == st_OFF) ? 1'b0 : 1'b1;

endmodule
// ****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.4 Simple FSM 2 (synchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_4.Simple_FSM_2_(synchronous reset)   // 無意義，快速找題目用
module top_module(
  input clk,
  input reset,    // synchronous reset to OFF
  input j,
  input k,
  output out
);

	parameter st_OFF=0;
  parameter st_ON=1;
  reg state;
  reg next_state;

  always @ (*) begin
  	if ( reset ) begin
  		 next_state = 0;
  	end else begin
  		case (state)
      st_OFF : next_state = (j) ? st_ON : st_OFF;
      st_ON  : next_state = (k) ? st_OFF: st_ON;
      default: next_state = (j) ? st_ON : st_OFF;
  		endcase

  	end
  end

  always @(posedge clk) begin
  	if ( reset ) begin
  		state <= st_OFF;
  	end else begin
  		state <= next_state;
  	end
  end

  assign out = (state == st_OFF) ? 1'b0 : 1'b1;

endmodule
// **********************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.5 Simple state transitions 3        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ********************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_5.Simple_state_transitions_3   // 無意義，快速找題目用
module top_module(
    input in,
    input [1:0] state,
    output [1:0] next_state,
    output out); //

    parameter A=0, B=1, C=2, D=3;

    // State transition logic: next_state = f(state, in)
    always @ (*) begin
    	case (state)
    		A : next_state = (in) ? B : A ;
    		B : next_state = (in) ? B : C ;
    		C : next_state = (in) ? D : A ;
    		D : next_state = (in) ? B : C ;
    		default : next_state = (in) ? B : A ;
    	endcase
    end

    // Output logic:  out = f(state) for a Moore state machine
    always @ (*) begin
    	case (state)
    		A : out = 0 ;
    		B : out = 0 ;
    		C : out = 0 ;
    		D : out = 1 ;
    		default : out = 0 ;
    	endcase
    end

endmodule

// ******************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.6 Simple one-hot state transitions 3        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_6 // 無意義，快速找題目用
module top_module(
    input in,
    input [3:0] state,
    output [3:0] next_state,
    output out); //

    parameter A=0;
    parameter B=1;
    parameter C=2;
    parameter D=3;

    // State transition logic: Derive an equation for each state flip-flop.
    assign next_state[A] =  (state[A] && ~in ) | (state[C] && ~in );
    assign next_state[B] =  (state[A] &&  in ) | (state[B] &&  in ) | (state[D] && in );
    assign next_state[C] =  (state[B] && ~in ) | (state[D] && ~in );
    assign next_state[D] =  (state[C] &&  in ) ;


    // Output logic:
    assign out = (state[D]) ? 1 : 0;

endmodule

// *****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.7 Simple FSM 3 (asynchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_7   // 無意義，快速找題目用
module top_module(
  input clk,
  input in,
  input areset,
  output out
); //

  reg [1:0] state;
  reg [1:0] next_state;

  parameter A=0, B=1, C=2, D=3;

  // State transition logic
  always @ (*) begin
  	if (areset) begin
  		next_state = A;
  	end else begin
  	  case (state)
    		A : next_state = (in) ? B : A ;
    		B : next_state = (in) ? B : C ;
    		C : next_state = (in) ? D : A ;
    		D : next_state = (in) ? B : C ;
    		default : next_state = A ;
  	  endcase

  	end
  end

  // State flip-flops with asynchronous reset
  always @(posedge clk or posedge areset) begin
	  if ( areset ) begin
	  	state <= A;
	  end else begin
	  	state <= next_state;
	  end
  end

  // Output logic
  always @ (*) begin
  	  case (state)
  	  	A : out = 0 ;
  	  	B : out = 0 ;
  	  	C : out = 0 ;
  	  	D : out = 1 ;
  	  	default : out = 0 ;
  	  endcase
  end

endmodule
// ****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.8 Simple FSM 3 (synchronous reset)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_8   // 無意義，快速找題目用
module top_module(
  input clk,
  input in,
  input reset,
  output out
); //

  reg [1:0] state;
  reg [1:0] next_state;

  parameter A=0, B=1, C=2, D=3;

  // State transition logic
  always @ (*) begin
  	 case (state)
    	A : next_state = (in) ? B : A ;
    	B : next_state = (in) ? B : C ;
    	C : next_state = (in) ? D : A ;
    	D : next_state = (in) ? B : C ;
    	default : next_state = A ;
  	 endcase
  end

  // State flip-flops with synchronous reset
  always @(posedge clk ) begin
	  if ( reset ) begin
	  	state <= A;
	  end else begin
	  	state <= next_state;
	  end
  end

  // Output logic
  always @ (*) begin
  	case (state)
  		A : out = 0 ;
  		B : out = 0 ;
  		C : out = 0 ;
  		D : out = 1 ;
  		default : out = 0 ;
  	endcase
  end

endmodule
// ***************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.9 Design a Moore FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
`define S03_2_5_9   // 無意義，快速找題目用
module top_module (
  input       clk,
  input       reset,
  input [3:1] s,
  output      fr3,
  output      fr2,
  output      fr1,
  output      dfr
);

parameter ST0 = 2'd0;
parameter ST1 = 2'd1;
parameter ST2 = 2'd2;
parameter ST3 = 2'd3;

reg [2:0] current;
reg [2:0] next_state;

always @ (*) begin
  case (current)
  	ST0 :
  	next_state = ( s == 3'b001 ) ? ST1 : ST0;
  	ST1 :
  	next_state = ( s == 3'b011) ? ST2 :
  	             ( s == 3'b000) ? ST0 : ST1;
  	ST2:
  	next_state = ( s == 3'b111) ? ST3 :
  	             ( s == 3'b001) ? ST1 : ST2;
  	ST3:
  	next_state = ( s == 3'b011) ? ST2 : ST3;

  	default : next_state = ST0;
  endcase
end

always @ (posedge clk ) begin
	if (reset) begin
		current <= ST0;
	end else begin
		current <= next_state;
	end
end


always @ (posedge clk ) begin
	if (reset) begin
    fr3 <= 1'b1;
    fr2 <= 1'b1;
    fr1 <= 1'b1;
    dfr <= 1'b1;
	end else begin
		case (next_state)
			ST0 : begin
				fr3 <= 1'b1;
        fr2 <= 1'b1;
        fr1 <= 1'b1;
        dfr <= 1'b1;
			end

			ST1 : begin
				fr3 <= 1'b0;
        fr2 <= 1'b1;
        fr1 <= 1'b1;
        dfr <= (current > next_state) ? 1'b1 :
               (current < next_state) ? 1'b0 : dfr;
			end

			ST2 : begin
				fr3 <= 1'b0;
        fr2 <= 1'b0;
        fr1 <= 1'b1;
        dfr <= (current > next_state) ? 1'b1 :
               (current < next_state) ? 1'b0 : dfr;
			end

			ST3 : begin
				fr3 <= 1'b0;
        fr2 <= 1'b0;
        fr1 <= 1'b0;
        dfr <= 1'b0;
			end


			default :  begin
				fr3 <= 1'b1;
        fr2 <= 1'b1;
        fr1 <= 1'b1;
        dfr <= 1'b1;
      end
		endcase

	end
end

endmodule
// *******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.10 Lemmings 1        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.11 Lemmings 2        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.12 Lemmings 3        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *******************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.13 Lemmings 4        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *****************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ********************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.14 One-hot FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ******************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ***************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.15 PS/2 packet parser        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ****************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.16 PS/2 packet parser and datapath        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.17 Serial receiver        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **********************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.18 Serial receiver and datapath        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***********************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *********************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.19 Serial receiver with parity checking        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *******************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *****************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.20 Sequence recognition        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *******************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.21 Q8: Design a Mealy FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *****************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ***************************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.22 Q5a: Serial two's complementer (Moore FSM)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *************************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ***************************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.23 Q5b: Serial two's complementer (Mealy FSM)        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *************************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *****************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.24 Q3a: FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *****************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.25 Q3b: FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ***********************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.26 Q3c: FSM logic        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// **********************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.27 Q6b: FSM next-state logic        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ********************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ******************************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.28 Q6c: FSM one-hot next-state logic        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ****************************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ****************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.29 Q6: FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// **************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *****************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.30 Q2a: FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// ***********************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.31 Q2b: One-hot FSM equations        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *****************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.32 Q2a: FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

// *************************************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//  S03-2-5.33 Q2b: Another FSM        /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// ***********************************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
